module HD(pc, clk, ONescrita, dadoEscrita, endereco, dadoLeitura, ck);
	input clk, ONescrita, ck;
	input [10:0] endereco, pc;
	input [31:0] dadoEscrita;
	output reg[31:0] dadoLeitura;
	reg [31:0] posHD	[1200:0];

	initial begin 
			/*KERNEL BLOCK*/


posHD[0] = 32'b00110100000000000000000000000001; /*jump    1  */
posHD[1] = 32'b00110100000000000000000000000010; /*JMP     2  */
posHD[2] = 32'b00100111100000000000000000000101;/*LOI    $28  5  */
posHD[3] = 32'b00001011100111000000000000000001;/*ADCI   $28 $28  1 */
posHD[4] = 32'b00100111010000000000000000000001;/*LOI    $26  1  */
posHD[5] = 32'b00100110000000000000000000000000;/*LOI    $16  0  */
posHD[6] = 32'b00100101000000000000000000000000;/*LOI    $8   0  */
posHD[7] = 32'b00100111001000000000000000110010;/*LOI    $25  50 */
posHD[8] = 32'b00100110111000000000000001000110;/*LOI    $23  70 */
posHD[9] = 32'b00100111000000000000000000000000;/*LOI    $24  0  */
posHD[10] = 32'b00100111011000000000000000000001;/*LOI    $27  1  */
posHD[11] = 32'b00100010111110101101100000000000; /*STWO   $23 $26  $27*/
posHD[12] = 32'b00100111110000000000001100100000;/*LOI    $30  800 */
posHD[13] = 32'b10011111011111100000000000000000;/*renameProgReg $27 $30  0 */
posHD[14] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[15] = 32'b00100111011000000000000000000010;/*LOI    $27  2  */
posHD[16] = 32'b00100010111110101101100000000000; /*STWO   $23 $26  $27*/
posHD[17] = 32'b00100111110000000000001101011100;/*LOI    $30  860 */
posHD[18] = 32'b10011111011111100000000000000000;/*renameProgReg $27 $30  0 */
posHD[19] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[20] = 32'b00100111011000000000000000000011;/*LOI    $27  3  */
posHD[21] = 32'b00100010111110101101100000000000; /*STWO   $23 $26  $27*/
posHD[22] = 32'b00100111110000000000001110011000;/*LOI    $30  920 */
posHD[23] = 32'b10011111011111100000000000000000;/*renameProgReg $27 $30  0 */
posHD[24] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[25] = 32'b00100111011000000000000000000100;/*LOI    $27  4  */
posHD[26] = 32'b00100010111110101101100000000000; /*STWO   $23 $26  $27*/
posHD[27] = 32'b00100111110000000000001111010100;/*LOI    $30  980 */
posHD[28] = 32'b10011111011111100000000000000000;/*renameProgReg $27 $30  0 */
posHD[29] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[30] = 32'b00100111011000000000000000000101;/*LOI    $27  5  */
posHD[31] = 32'b00100010111110101101100000000000; /*STWO   $23 $26  $27*/
posHD[32] = 32'b00100111110000000000010000010000;/*LOI    $30  1040 */
posHD[33] = 32'b10011111011111100000000000000000;/*renameProgReg $27 $30  0 */
posHD[34] = 32'b10001000000000000000000000001011; /*li6     11 */
posHD[35] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[36] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[37] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[38] = 32'b01000011110111110000000000101011;/*BNEQ   $30 $31  43*/
posHD[39] = 32'b10001000000000000000000000001101; /*li6     13 */
posHD[40] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[41] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[42] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[43] = 32'b00100111110000000000000000000010;/*LOI    $30  2  */
posHD[44] = 32'b01000011110111110000000000110001;/*BNEQ   $30 $31  49*/
posHD[45] = 32'b10001000000000000000000000001110; /*li6     14 */
posHD[46] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[47] = 32'b00110100000000000000000001110010; /*JMP     114 */
posHD[48] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[49] = 32'b00100111110000000000000000000011;/*LOI    $30  3  */
posHD[50] = 32'b01000011110111110000000000110111;/*BNEQ   $30 $31  55*/
posHD[51] = 32'b10001000000000000000000000001111; /*li6     15 */
posHD[52] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[53] = 32'b00110100000000000000000000111101; /*JMP     61 */
posHD[54] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[55] = 32'b00100111110000000000000000000100;/*LOI    $30  4  */
posHD[56] = 32'b01000011110111110000000000100010;/*BNEQ   $30 $31  34*/
posHD[57] = 32'b10001000000000000000000000010000; /*li6     16 */
posHD[58] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[59] = 32'b00110100000000000000000001011111; /*JMP     95 */
posHD[60] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[61] = 32'b10001000000000000000000000010011; /*li6     19 */
posHD[62] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[63] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[64] = 32'b00100111010000000000000000000001;/*LOI    $26  1  */
posHD[65] = 32'b01001011010111001110100000000000; /*SLET   $26 $28  $29*/
posHD[66] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[67] = 32'b01000011101111100000000001011101;/*BNEQ   $29 $30  93*/
posHD[68] = 32'b00011110111110101111000000000000; /*LOWO   $23 $26  $30*/
posHD[69] = 32'b01000011111111100000000001011011;/*BNEQ   $31 $30  91*/
posHD[70] = 32'b10011011110101010000000000000000;/*switchCtx $30 $21  0 */
posHD[71] = 32'b00101011110110110000000000000000;/*MOV    $30 $27  0 */
posHD[72] = 32'b10001000000000000000000000010100; /*li6     20 */
posHD[73] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[74] = 32'b01010010100000000000000000000000;/*IN     $20  0  */
posHD[75] = 32'b00100100011000000000000000000001;/*LOI    $3   1  */
posHD[76] = 32'b01001000011111001110100000000000; /*SLET   $3  $28  $29*/
posHD[77] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[78] = 32'b01000011101111100000000001010110;/*BNEQ   $29 $30  86*/
posHD[79] = 32'b00011110111000111111000000000000; /*LOWO   $23 $3   $30*/
posHD[80] = 32'b01000010100111100000000001010100;/*BNEQ   $20 $30  84*/
posHD[81] = 32'b10001000000000000000000000011010; /*li6     26 */
posHD[82] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[83] = 32'b00110100000000000000000001001010; /*JMP     74 */
posHD[84] = 32'b00001000011000110000000000000001;/*ADCI   $3  $3   1 */
posHD[85] = 32'b00110100000000000000000001001100; /*JMP     76 */
posHD[86] = 32'b10011110100101010000000000000000;/*renameProgReg $20 $21  0 */
posHD[87] = 32'b00100010111110101010000000000000; /*STWO   $23 $26  $20*/
posHD[88] = 32'b10001000000000000000000000010100; /*li6     20 */
posHD[89] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[90] = 32'b00110100000000000000000001011100; /*JMP     92 */
posHD[91] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[92] = 32'b00110100000000000000000001000001; /*JMP     65 */
posHD[93] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[94] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[95] = 32'b10001000000000000000000000010101; /*li6     21 */
posHD[96] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[97] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[98] = 32'b00101011111101000000000000000000;/*MOV    $31 $20  0 */
posHD[99] = 32'b00100111010000000000000000000001;/*LOI    $26  1  */
posHD[100] = 32'b01001011010111001110100000000000; /*SLET   $26 $28  $29*/
posHD[101] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[102] = 32'b01000011101111100000000001110000;/*BNEQ   $29 $30  112*/
posHD[103] = 32'b00011110111110101111000000000000; /*LOWO   $23 $26  $30*/
posHD[104] = 32'b01000011111111100000000001101110;/*BNEQ   $31 $30  110*/
posHD[105] = 32'b10001000000000000000000000010110; /*li6     22 */
posHD[106] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[107] = 32'b00100111110000000000000000000000;/*LOI    $30  0  */
posHD[108] = 32'b00100010111110101111000000000000; /*STWO   $23 $26  $30*/
posHD[109] = 32'b00110100000000000000000001110000; /*JMP     112 */
posHD[110] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[111] = 32'b00110100000000000000000001100100; /*JMP     100 */
posHD[112] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[113] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[114] = 32'b10001000000000000000000000011011; /*li6     27 */
posHD[115] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[116] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[117] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[118] = 32'b00100111101000000000000000000010;/*LOI    $29  2  */
posHD[119] = 32'b01000011111111100000000011111001;/*BNEQ   $31 $30  249*/
posHD[120] = 32'b10001000000000000000000000011100; /*li6     28 */
posHD[121] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[122] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[123] = 32'b00100111010000000000000000000001;/*LOI    $26  1  */
posHD[124] = 32'b01001011010111001111000000000000; /*SLET   $26 $28  $30*/
posHD[125] = 32'b00100111101000000000000000000001;/*LOI    $29  1  */
posHD[126] = 32'b01000011101111100000000000100010;/*BNEQ   $29 $30  34*/
posHD[127] = 32'b00011110111110101101100000000000; /*LOWO   $23 $26  $27*/
posHD[128] = 32'b01000011111110110000000011110111;/*BNEQ   $31 $27  247*/
posHD[129] = 32'b10011011011101010000000000000000;/*switchCtx $27 $21  0 */
posHD[130] = 32'b01110010101000000000001111101000; /*COPY    21, 1000*/
posHD[131] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[132] = 32'b01110010101000000000001111101001; /*COPY    21, 1001*/
posHD[133] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[134] = 32'b01110010101000000000001111101010; /*COPY    21, 1002*/
posHD[135] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[136] = 32'b01110010101000000000001111101011; /*COPY    21, 1003*/
posHD[137] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[138] = 32'b01110010101000000000001111101100; /*COPY    21, 1004*/
posHD[139] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[140] = 32'b01110010101000000000001111101101; /*COPY    21, 1005*/
posHD[141] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[142] = 32'b01110010101000000000001111101110; /*COPY    21, 1006*/
posHD[143] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[144] = 32'b01110010101000000000001111101111; /*COPY    21, 1007*/
posHD[145] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[146] = 32'b01110010101000000000001111110000; /*COPY    21, 1008*/
posHD[147] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[148] = 32'b01110010101000000000001111110001; /*COPY    21, 1009*/
posHD[149] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[150] = 32'b01110010101000000000001111110010; /*COPY    21, 1010*/
posHD[151] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[152] = 32'b01110010101000000000001111110011; /*COPY    21, 1011*/
posHD[153] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[154] = 32'b01110010101000000000001111110100; /*COPY    21, 1012*/
posHD[155] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[156] = 32'b01110010101000000000001111110101; /*COPY    21, 1013*/
posHD[157] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[158] = 32'b01110010101000000000001111110110; /*COPY    21, 1014*/
posHD[159] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[160] = 32'b01110010101000000000001111110111; /*COPY    21, 1015*/
posHD[161] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[162] = 32'b01110010101000000000001111111000; /*COPY    21, 1016*/
posHD[163] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[164] = 32'b01110010101000000000001111111001; /*COPY    21, 1017*/
posHD[165] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[166] = 32'b01110010101000000000001111111010; /*COPY    21, 1018*/
posHD[167] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[168] = 32'b01110010101000000000001111111011; /*COPY    21, 1019*/
posHD[169] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[170] = 32'b01110010101000000000001111111100; /*COPY    21, 1020*/
posHD[171] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[172] = 32'b01110010101000000000001111111101; /*COPY    21, 1021*/
posHD[173] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[174] = 32'b01110010101000000000001111111110; /*COPY    21, 1022*/
posHD[175] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[176] = 32'b01110010101000000000001111111111; /*COPY    21, 1023*/
posHD[177] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[178] = 32'b01110010101000000000010000000000; /*COPY    21, 1024*/
posHD[179] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[180] = 32'b01110010101000000000010000000001; /*COPY    21, 1025*/
posHD[181] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[182] = 32'b01110010101000000000010000000010; /*COPY    21, 1026*/
posHD[183] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[184] = 32'b01110010101000000000010000000011; /*COPY    21, 1027*/
posHD[185] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[186] = 32'b01110010101000000000010000000100; /*COPY    21, 1028*/
posHD[187] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[188] = 32'b01110010101000000000010000000101; /*COPY    21, 1029*/
posHD[189] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[190] = 32'b01110010101000000000010000000110; /*COPY    21, 1030*/
posHD[191] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[192] = 32'b01110010101000000000010000000111; /*COPY    21, 1031*/
posHD[193] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[194] = 32'b01110010101000000000010000001000; /*COPY    21, 1032*/
posHD[195] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[196] = 32'b01110010101000000000010000001001; /*COPY    21, 1033*/
posHD[197] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[198] = 32'b01110010101000000000010000001010; /*COPY    21, 1034*/
posHD[199] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[200] = 32'b01110010101000000000010000001011; /*COPY    21, 1035*/
posHD[201] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[202] = 32'b01110010101000000000010000001100; /*COPY    21, 1036*/
posHD[203] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[204] = 32'b01110010101000000000010000001101; /*COPY    21, 1037*/
posHD[205] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[206] = 32'b01110010101000000000010000001110; /*COPY    21, 1038*/
posHD[207] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[208] = 32'b01110010101000000000010000001111; /*COPY    21, 1039*/
posHD[209] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[210] = 32'b01110010101000000000010000010000; /*COPY    21, 1040*/
posHD[211] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[212] = 32'b01110010101000000000010000010001; /*COPY    21, 1041*/
posHD[213] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[214] = 32'b01110010101000000000010000010010; /*COPY    21, 1042*/
posHD[215] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[216] = 32'b01110010101000000000010000010011; /*COPY    21, 1043*/
posHD[217] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[218] = 32'b01110010101000000000010000010100; /*COPY    21, 1044*/
posHD[219] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[220] = 32'b01110010101000000000010000010101; /*COPY    21, 1045*/
posHD[221] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[222] = 32'b01110010101000000000010000010110; /*COPY    21, 1046*/
posHD[223] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[224] = 32'b01110010101000000000010000010111; /*COPY    21, 1047*/
posHD[225] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[226] = 32'b01110010101000000000010000011000; /*COPY    21, 1048*/
posHD[227] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[228] = 32'b01110010101000000000010000011001; /*COPY    21, 1049*/
posHD[229] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[230] = 32'b01110010101000000000010000011010; /*COPY    21, 1050*/
posHD[231] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[232] = 32'b01110010101000000000010000011011; /*COPY    21, 1051*/
posHD[233] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[234] = 32'b01110010101000000000010000011100; /*COPY    21, 1052*/
posHD[235] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[236] = 32'b01110010101000000000010000011101; /*COPY    21, 1053*/
posHD[237] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[238] = 32'b01110010101000000000010000011110; /*COPY    21, 1054*/
posHD[239] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[240] = 32'b01110010101000000000010000011111; /*COPY    21, 1055*/
posHD[241] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[242] = 32'b01110010101000000000010000100000; /*COPY    21, 1056*/
posHD[243] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[244] = 32'b00100110101000000000010001001100;/*LOI    $21  1100 */
posHD[245] = 32'b01110010101000000000010000100001; /*COPY    21, 1057*/
posHD[246] = 32'b00110100000000000000001111101000; /*JMP     1000 */
posHD[247] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[248] = 32'b00110100000000000000000001111100; /*JMP     124 */
posHD[249] = 32'b10001000000000000000000000010001; /*li6     17 */
posHD[250] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[251] = 32'b00100110100000000000000000000000;/*LOI    $20  0  */
posHD[252] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[253] = 32'b00101011111101100000000000000000;/*MOV    $31 $22  0 */
posHD[254] = 32'b00100100111000000000000000000000;/*LOI    $7   0  */
posHD[255] = 32'b01001000111101101110100000000000; /*SLET   $7  $22  $29*/
posHD[256] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[257] = 32'b01000011101111100000000100010001;/*BNEQ   $29 $30  273*/
posHD[258] = 32'b10001000000000000000000000010010; /*li6     18 */
posHD[259] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[260] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[261] = 32'b00100111010000000000000000000001;/*LOI    $26  1  */
posHD[262] = 32'b01001011010111001111000000000000; /*SLET   $26 $28  $30*/
posHD[263] = 32'b00100111101000000000000000000001;/*LOI    $29  1  */
posHD[264] = 32'b01000011101111100000000011111111;/*BNEQ   $29 $30  255*/
posHD[265] = 32'b00011110111110101111000000000000; /*LOWO   $23 $26  $30*/
posHD[266] = 32'b01000011110111110000000100001101;/*BNEQ   $30 $31  269*/
posHD[267] = 32'b00100011001001111111100000000000; /*STWO   $25 $7   $31*/
posHD[268] = 32'b00110100000000000000000100001111; /*JMP     271 */
posHD[269] = 32'b00001011010110100000000000000001;/*ADCI   $26 $26  1 */
posHD[270] = 32'b00110100000000000000000100000110; /*JMP     262 */
posHD[271] = 32'b00001000111001110000000000000001;/*ADCI   $7  $7   1 */
posHD[272] = 32'b00110100000000000000000011111111; /*JMP     255 */
posHD[273] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[274] = 32'b10001000000000000000000000010111; /*li6     23 */
posHD[275] = 32'b10000100000000000000000000000000; /*emit    0  */
posHD[276] = 32'b00100100111000000000000000000000;/*LOI    $7   0  */
posHD[277] = 32'b01001000111101101111000000000000; /*SLET   $7  $22  $30*/
posHD[278] = 32'b00100111101000000000000000000001;/*LOI    $29  1  */
posHD[279] = 32'b01000011101111100000000111000000;/*BNEQ   $29 $30  448*/
posHD[280] = 32'b00011111001001111111000000000000; /*LOWO   $25 $7   $30*/
posHD[281] = 32'b00101011110110110000000000000000;/*MOV    $30 $27  0 */
posHD[282] = 32'b01010111011000000000000000000000;/*OUT    $27  0  */
posHD[283] = 32'b10011011011101010000000000000000;/*switchCtx $27 $21  0 */
posHD[284] = 32'b01110010101000000000001111101000; /*COPY    21, 1000*/
posHD[285] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[286] = 32'b01110010101000000000001111101001; /*COPY    21, 1001*/
posHD[287] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[288] = 32'b01110010101000000000001111101010; /*COPY    21, 1002*/
posHD[289] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[290] = 32'b01110010101000000000001111101011; /*COPY    21, 1003*/
posHD[291] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[292] = 32'b01110010101000000000001111101100; /*COPY    21, 1004*/
posHD[293] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[294] = 32'b01110010101000000000001111101101; /*COPY    21, 1005*/
posHD[295] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[296] = 32'b01110010101000000000001111101110; /*COPY    21, 1006*/
posHD[297] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[298] = 32'b01110010101000000000001111101111; /*COPY    21, 1007*/
posHD[299] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[300] = 32'b01110010101000000000001111110000; /*COPY    21, 1008*/
posHD[301] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[302] = 32'b01110010101000000000001111110001; /*COPY    21, 1009*/
posHD[303] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[304] = 32'b01110010101000000000001111110010; /*COPY    21, 1010*/
posHD[305] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[306] = 32'b01110010101000000000001111110011; /*COPY    21, 1011*/
posHD[307] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[308] = 32'b01110010101000000000001111110100; /*COPY    21, 1012*/
posHD[309] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[310] = 32'b01110010101000000000001111110101; /*COPY    21, 1013*/
posHD[311] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[312] = 32'b01110010101000000000001111110110; /*COPY    21, 1014*/
posHD[313] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[314] = 32'b01110010101000000000001111110111; /*COPY    21, 1015*/
posHD[315] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[316] = 32'b01110010101000000000001111111000; /*COPY    21, 1016*/
posHD[317] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[318] = 32'b01110010101000000000001111111001; /*COPY    21, 1017*/
posHD[319] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[320] = 32'b01110010101000000000001111111010; /*COPY    21, 1018*/
posHD[321] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[322] = 32'b01110010101000000000001111111011; /*COPY    21, 1019*/
posHD[323] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[324] = 32'b01110010101000000000001111111100; /*COPY    21, 1020*/
posHD[325] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[326] = 32'b01110010101000000000001111111101; /*COPY    21, 1021*/
posHD[327] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[328] = 32'b01110010101000000000001111111110; /*COPY    21, 1022*/
posHD[329] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[330] = 32'b01110010101000000000001111111111; /*COPY    21, 1023*/
posHD[331] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[332] = 32'b01110010101000000000010000000000; /*COPY    21, 1024*/
posHD[333] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[334] = 32'b01110010101000000000010000000001; /*COPY    21, 1025*/
posHD[335] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[336] = 32'b01110010101000000000010000000010; /*COPY    21, 1026*/
posHD[337] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[338] = 32'b01110010101000000000010000000011; /*COPY    21, 1027*/
posHD[339] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[340] = 32'b01110010101000000000010000000100; /*COPY    21, 1028*/
posHD[341] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[342] = 32'b01110010101000000000010000000101; /*COPY    21, 1029*/
posHD[343] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[344] = 32'b01110010101000000000010000000110; /*COPY    21, 1030*/
posHD[345] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[346] = 32'b01110010101000000000010000000111; /*COPY    21, 1031*/
posHD[347] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[348] = 32'b01110010101000000000010000001000; /*COPY    21, 1032*/
posHD[349] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[350] = 32'b01110010101000000000010000001001; /*COPY    21, 1033*/
posHD[351] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[352] = 32'b01110010101000000000010000001010; /*COPY    21, 1034*/
posHD[353] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[354] = 32'b01110010101000000000010000001011; /*COPY    21, 1035*/
posHD[355] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[356] = 32'b01110010101000000000010000001100; /*COPY    21, 1036*/
posHD[357] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[358] = 32'b01110010101000000000010000001101; /*COPY    21, 1037*/
posHD[359] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[360] = 32'b01110010101000000000010000001110; /*COPY    21, 1038*/
posHD[361] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[362] = 32'b01110010101000000000010000001111; /*COPY    21, 1039*/
posHD[363] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[364] = 32'b01110010101000000000010000010000; /*COPY    21, 1040*/
posHD[365] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[366] = 32'b01110010101000000000010000010001; /*COPY    21, 1041*/
posHD[367] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[368] = 32'b01110010101000000000010000010010; /*COPY    21, 1042*/
posHD[369] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[370] = 32'b01110010101000000000010000010011; /*COPY    21, 1043*/
posHD[371] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[372] = 32'b01110010101000000000010000010100; /*COPY    21, 1044*/
posHD[373] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[374] = 32'b01110010101000000000010000010101; /*COPY    21, 1045*/
posHD[375] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[376] = 32'b01110010101000000000010000010110; /*COPY    21, 1046*/
posHD[377] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[378] = 32'b01110010101000000000010000010111; /*COPY    21, 1047*/
posHD[379] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[380] = 32'b01110010101000000000010000011000; /*COPY    21, 1048*/
posHD[381] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[382] = 32'b01110010101000000000010000011001; /*COPY    21, 1049*/
posHD[383] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[384] = 32'b01110010101000000000010000011010; /*COPY    21, 1050*/
posHD[385] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[386] = 32'b01110010101000000000010000011011; /*COPY    21, 1051*/
posHD[387] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[388] = 32'b01110010101000000000010000011100; /*COPY    21, 1052*/
posHD[389] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[390] = 32'b01110010101000000000010000011101; /*COPY    21, 1053*/
posHD[391] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[392] = 32'b01110010101000000000010000011110; /*COPY    21, 1054*/
posHD[393] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[394] = 32'b01110010101000000000010000011111; /*COPY    21, 1055*/
posHD[395] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[396] = 32'b01110010101000000000010000100000; /*COPY    21, 1056*/
posHD[397] = 32'b00001010101101010000000000000001;/*ADCI   $21 $21  1 */
posHD[398] = 32'b01110100111000000000000000000000;/*LR     $7   0  */
posHD[399] = 32'b01110100111000000000000000000001;/*LR     $7   1  */
posHD[400] = 32'b01110100111000000000000000000010;/*LR     $7   2  */
posHD[401] = 32'b01110100111000000000000000000011;/*LR     $7   3  */
posHD[402] = 32'b01110100111000000000000000000100;/*LR     $7   4  */
posHD[403] = 32'b01110100111000000000000000000101;/*LR     $7   5  */
posHD[404] = 32'b01110100111000000000000000000110;/*LR     $7   6  */
posHD[405] = 32'b01110100111000000000000000001000;/*LR     $7   8  */
posHD[406] = 32'b01110100111000000000000000001001;/*LR     $7   9  */
posHD[407] = 32'b01110100111000000000000000001010;/*LR     $7   10 */
posHD[408] = 32'b01110100111000000000000000001011;/*LR     $7   11 */
posHD[409] = 32'b01110100111000000000000000001100;/*LR     $7   12 */
posHD[410] = 32'b01110100111000000000000000001101;/*LR     $7   13 */
posHD[411] = 32'b01110100111000000000000000001110;/*LR     $7   14 */
posHD[412] = 32'b01110100111000000000000000001111;/*LR     $7   15 */
posHD[413] = 32'b01110100111000000000000000010001;/*LR     $7   17 */
posHD[414] = 32'b01110100111000000000000000010010;/*LR     $7   18 */
posHD[415] = 32'b01110100111000000000000000010011;/*LR     $7   19 */
posHD[416] = 32'b01110100111000000000000000011101;/*LR     $7   29 */
posHD[417] = 32'b01110100111000000000000000011110;/*LR     $7   30 */
posHD[418] = 32'b01110100111000000000000000011111;/*LR     $7   31 */
posHD[419] = 32'b00100111110000000000000000000000;/*LOI    $30  0  */
posHD[420] = 32'b01000011110100000000000110100111;/*BNEQ   $30 $16  423*/
posHD[421] = 32'b00100101000000000000000000000000;/*LOI    $8   0  */
posHD[422] = 32'b00001001000010000000001111100111;/*ADCI   $8  $8   999*/
posHD[423] = 32'b00011000000000000000000000000000; /*CPC     0  */
posHD[424] = 32'b00111001000000000000000000000000;/*JMPR   $8   0  */
posHD[425] = 32'b01111000111000000000000000000000;/*SR     $7   0  */
posHD[426] = 32'b01111000111000000000000000000001;/*SR     $7   1  */
posHD[427] = 32'b01111000111000000000000000000010;/*SR     $7   2  */
posHD[428] = 32'b01111000111000000000000000000011;/*SR     $7   3  */
posHD[429] = 32'b01111000111000000000000000000100;/*SR     $7   4  */
posHD[430] = 32'b01111000111000000000000000000101;/*SR     $7   5  */
posHD[431] = 32'b01111000111000000000000000000110;/*SR     $7   6  */
posHD[432] = 32'b01111000111000000000000000001000;/*SR     $7   8  */
posHD[433] = 32'b01111000111000000000000000001001;/*SR     $7   9  */
posHD[434] = 32'b01111000111000000000000000001010;/*SR     $7   10 */
posHD[435] = 32'b01111000111000000000000000001011;/*SR     $7   11 */
posHD[436] = 32'b01111000111000000000000000001100;/*SR     $7   12 */
posHD[437] = 32'b01111000111000000000000000001101;/*SR     $7   13 */
posHD[438] = 32'b01111000111000000000000000001110;/*SR     $7   14 */
posHD[439] = 32'b01111000111000000000000000001111;/*SR     $7   15 */
posHD[440] = 32'b01111000111000000000000000010001;/*SR     $7   17 */
posHD[441] = 32'b01111000111000000000000000010010;/*SR     $7   18 */
posHD[442] = 32'b01111000111000000000000000010011;/*SR     $7   19 */
posHD[443] = 32'b01111000111000000000000000011101;/*SR     $7   29 */
posHD[444] = 32'b01111000111000000000000000011110;/*SR     $7   30 */
posHD[445] = 32'b01111000111000000000000000011111;/*SR     $7   31 */
posHD[446] = 32'b00001000111001110000000000000001;/*ADCI   $7  $7   1 */
posHD[447] = 32'b00110100000000000000000100010101; /*JMP     277 */
posHD[448] = 32'b00100110000000000000000000001010;/*LOI    $16  10 */
posHD[449] = 32'b00100100111000000000000000000000;/*LOI    $7   0  */
posHD[450] = 32'b00110100000000000000000100010101; /*JMP     277 */
posHD[451] = 32'b01011100000000000000000000000000; /*HALT    0  */
posHD[452] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[453] = 32'b00100111000000000000000000000000;/*LOI    $24  0  */
posHD[454] = 32'b00001011000110000000000000000001;/*ADCI   $24 $24  1 */
posHD[455] = 32'b00110100000000000000000110111110; /*JMP     446 */
posHD[456] = 32'b00110100000000000000000111000100; /*JMP     452 */
posHD[457] = 32'b01011100000000000000000000000000; /*HALT    0  */

  
		/*SAVED BLOCK*/


		/*INSTRUCTION BLOCK*/
//fatorial

posHD[800] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[801] = 32'b00110100000000000000010000000011; /*JMP    $1027*/
posHD[802] = 32'b00100101001000000000000000000001;/*LOI    $9   1  */
posHD[803] = 32'b00101000000111100000000000000000;/*MOV    $0  $30  0 */
posHD[804] = 32'b00101000100100010000000000000000;/*MOV    $4  $17  0 */
posHD[805] = 32'b00101000100111010000000000000000;/*MOV    $4  $29  0 */
posHD[806] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[807] = 32'b00100111110000000000000000000000;/*LOI    $30  0  */
posHD[808] = 32'b01001111101111101110100000000000; /*SGRT   $29 $30  $29*/
posHD[809] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[810] = 32'b01000011110111010000001111111110;/*BNEQ   $30 $29  1022*/
posHD[811] = 32'b00101001001100010000000000000000;/*MOV    $9  $17  0 */
posHD[812] = 32'b00101000100111010000000000000000;/*MOV    $4  $29  0 */
posHD[813] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[814] = 32'b01100011101111101111000000000000; /*MULT   $29 $30  $30*/
posHD[815] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[816] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[817] = 32'b00101000100100010000000000000000;/*MOV    $4  $17  0 */
posHD[818] = 32'b00101010001111010000000000000000;/*MOV    $17 $29  0 */
posHD[819] = 32'b00001111101111100000000000000001;/*SUBI   $29 $30  1 */
posHD[820] = 32'b00101011110001000000000000000000;/*MOV    $30 $4   0 */
posHD[821] = 32'b00110100000000000000001111101100; /*JMP     1004 */
posHD[822] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[823] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[824] = 32'b00101001001111110000000000000000;/*MOV    $9  $31  0 */
posHD[825] = 32'b01010111111000000000000000000000;/*OUT    $31  0  */
posHD[826] = 32'b00111000000000000000000000000000;/*JMPR   $0   0  */
posHD[827] = 32'b00110100000000000000010000000100; /*JMP     1028 */
posHD[828] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[829] = 32'b00101000000111100000000000000000;/*MOV    $0  $30  0 */
posHD[830] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[831] = 32'b00101011110000000000000000000000;/*MOV    $30 $0   0 */
posHD[832] = 32'b00101000000001000000000000000000;/*MOV    $0  $4   0 */
posHD[833] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[834] = 32'b01101000000000000000001111101010; /*JAL     1002 */
posHD[835] = 32'b00101000000111110000000000000000;/*MOV    $0  $31  0 */
posHD[836] = 32'b10100000000000000000000000000000; /*interrupCPC     0  */


//gcd

posHD[860] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[861] = 32'b00110100000000000000010000000011; /*JMP    $1027*/
posHD[862] = 32'b00101000101100010000000000000000;/*MOV    $5  $17  0 */
posHD[863] = 32'b00101000101111010000000000000000;/*MOV    $5  $29  0 */
posHD[864] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[865] = 32'b00100111101000000000000000000000;/*LOI    $29  0  */
posHD[866] = 32'b01000011110111010000001111110001;/*BNEQ   $30 $29  1009*/
posHD[867] = 32'b00101000100000010000000000000000;/*MOV    $4  $1   0 */
posHD[868] = 32'b00110100000000000000010000000001; /*JMP     1025 */
posHD[869] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[870] = 32'b00101000100111100000000000000000;/*MOV    $4  $30  0 */
posHD[871] = 32'b00101000101001000000000000000000;/*MOV    $5  $4   0 */
posHD[872] = 32'b00101011110011110000000000000000;/*MOV    $30 $15  0 */
posHD[873] = 32'b00101001111100010000000000000000;/*MOV    $15 $17  0 */
posHD[874] = 32'b00101001111100100000000000000000;/*MOV    $15 $18  0 */
posHD[875] = 32'b00101000101111010000000000000000;/*MOV    $5  $29  0 */
posHD[876] = 32'b00101010010111100000000000000000;/*MOV    $18 $30  0 */
posHD[877] = 32'b01101111110111011111000000000000; /*DIV    $30 $29  $30*/
posHD[878] = 32'b00101000101100100000000000000000;/*MOV    $5  $18  0 */
posHD[879] = 32'b00101010010111010000000000000000;/*MOV    $18 $29  0 */
posHD[880] = 32'b01100011101111101111000000000000; /*MULT   $29 $30  $30*/
posHD[881] = 32'b00101010001111010000000000000000;/*MOV    $17 $29  0 */
posHD[882] = 32'b00000111101111101111000000000000; /*SUB    $29 $30  $30*/
posHD[883] = 32'b00101011110001010000000000000000;/*MOV    $30 $5   0 */
posHD[884] = 32'b00110100000000000000001111101010; /*JMP     1002 */
posHD[885] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[886] = 32'b00111000000000000000000000000000;/*JMPR   $0   0  */
posHD[887] = 32'b00110100000000000000010000000100; /*JMP     1028 */
posHD[888] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[889] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[890] = 32'b00101001001111100000000000000000;/*MOV    $9  $30  0 */
posHD[891] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[892] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[893] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[894] = 32'b00101001001111100000000000000000;/*MOV    $9  $30  0 */
posHD[895] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[896] = 32'b00101011110010100000000000000000;/*MOV    $30 $10  0 */
posHD[897] = 32'b00101001001111110000000000000000;/*MOV    $9  $31  0 */
posHD[898] = 32'b00101001001001000000000000000000;/*MOV    $9  $4   0 */
posHD[899] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[900] = 32'b00101001010111110000000000000000;/*MOV    $10 $31  0 */
posHD[901] = 32'b00101011111010100000000000000000;/*MOV    $31 $10  0 */
posHD[902] = 32'b00101001010001010000000000000000;/*MOV    $10 $5   0 */
posHD[903] = 32'b01101000000000000000001111101010; /*JAL     1002 */
posHD[904] = 32'b00101000001111110000000000000000;/*MOV    $1  $31  0 */
posHD[905] = 32'b01010111111000000000000000000000;/*OUT    $31  0  */

posHD[906] = 32'b10100000000000000000000000000000; /*interrupCPC     0  */



//somaVet
posHD[920] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[921] = 32'b00110100000000000000010000000101; /*JMP    $1029*/
posHD[922] = 32'b00100101010000000000000000000000;/*LOI    $10  0  */
posHD[923] = 32'b00101000000111100000000000000000;/*MOV    $0  $30  0 */
posHD[924] = 32'b00100101001000000000000000000000;/*LOI    $9   0  */
posHD[925] = 32'b00101001001111100000000000000000;/*MOV    $9  $30  0 */
posHD[926] = 32'b00101001001100010000000000000000;/*MOV    $9  $17  0 */
posHD[927] = 32'b00101001001111010000000000000000;/*MOV    $9  $29  0 */
posHD[928] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[929] = 32'b00100111110000000000000000000100;/*LOI    $30  4  */
posHD[930] = 32'b01001011101111101110100000000000; /*SLET   $29 $30  $29*/
posHD[931] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[932] = 32'b01000011110111010000010000000010;/*BNEQ   $30 $29  1026*/
posHD[933] = 32'b00011100100010011110100000000000; /*LOWO   $4  $9   $29*/
posHD[934] = 32'b00101001001100100000000000000000;/*MOV    $9  $18  0 */
posHD[935] = 32'b00101001001111100000000000000000;/*MOV    $9  $30  0 */
posHD[936] = 32'b00101001010111100000000000000000;/*MOV    $10 $30  0 */
posHD[937] = 32'b00000011101111101111000000000000; /*ADC    $29 $30  $30*/
posHD[938] = 32'b00101011110010100000000000000000;/*MOV    $30 $10  0 */
posHD[939] = 32'b00101011110010100000000000000000;/*MOV    $30 $10  0 */
posHD[940] = 32'b00101001001100110000000000000000;/*MOV    $9  $19  0 */
posHD[941] = 32'b00101010011111010000000000000000;/*MOV    $19 $29  0 */
posHD[942] = 32'b00001011101111100000000000000001;/*ADCI   $29 $30  1 */
posHD[943] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[944] = 32'b00110100000000000000001111101110; /*JMP     1006 */
posHD[945] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[946] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[947] = 32'b00101001010000010000000000000000;/*MOV    $10 $1   0 */
posHD[948] = 32'b00111000000000000000000000000000;/*JMPR   $0   0  */
posHD[949] = 32'b00110100000000000000010000000110; /*JMP     1030 */
posHD[950] = 32'b00100100001000000000000000000000;/*LOI    $1   0  */
posHD[951] = 32'b00101000001111100000000000000000;/*MOV    $1  $30  0 */
posHD[952] = 32'b00101000001100010000000000000000;/*MOV    $1  $17  0 */
posHD[953] = 32'b00101000001111010000000000000000;/*MOV    $1  $29  0 */
posHD[954] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[955] = 32'b00100111110000000000000000000100;/*LOI    $30  4  */
posHD[956] = 32'b01001011101111101110100000000000; /*SLET   $29 $30  $29*/
posHD[957] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[958] = 32'b01000011110111010000010000011010;/*BNEQ   $30 $29  1050*/
posHD[959] = 32'b00011100010000011111000000000000; /*LOWO   $2  $1   $30*/
posHD[960] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[961] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[962] = 32'b00100000010000011111000000000000; /*STWO   $2  $1   $30*/
posHD[963] = 32'b00101000001100010000000000000000;/*MOV    $1  $17  0 */
posHD[964] = 32'b00101000001111010000000000000000;/*MOV    $1  $29  0 */
posHD[965] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[966] = 32'b00001011101111100000000000000001;/*ADCI   $29 $30  1 */
posHD[967] = 32'b00101011110000010000000000000000;/*MOV    $30 $1   0 */
posHD[968] = 32'b00110100000000000000010000001000; /*JMP     1032 */
posHD[969] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[970] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[971] = 32'b00101000010111110000000000000000;/*MOV    $2  $31  0 */
posHD[972] = 32'b00101000010001000000000000000000;/*MOV    $2  $4   0 */
posHD[973] = 32'b01101000000000000000001111101010; /*JAL     1002 */
posHD[974] = 32'b00101000001111110000000000000000;/*MOV    $1  $31  0 */
posHD[975] = 32'b01010111111000000000000000000000;/*OUT    $31  0  */
posHD[976] = 32'b10100000000000000000000000000000; /*interrupCPC     0  */


//media
posHD[980] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[981] = 32'b00110100000000000000001111111000; /*JMP    $1016*/
posHD[982] = 32'b00101000100100010000000000000000;/*MOV    $4  $17  0 */
posHD[983] = 32'b00101000101111010000000000000000;/*MOV    $5  $29  0 */
posHD[984] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[985] = 32'b00000011101111101111000000000000; /*ADC    $29 $30  $30*/
posHD[986] = 32'b00101011110010100000000000000000;/*MOV    $30 $10  0 */
posHD[987] = 32'b00101011110010100000000000000000;/*MOV    $30 $10  0 */
posHD[988] = 32'b00101001010100010000000000000000;/*MOV    $10 $17  0 */
posHD[989] = 32'b00101010001111010000000000000000;/*MOV    $17 $29  0 */
posHD[990] = 32'b00100111110000000000000000000010;/*LOI    $30  2  */
posHD[991] = 32'b01101111101111101111000000000000; /*DIV    $29 $30  $30*/
posHD[992] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[993] = 32'b00101001001111110000000000000000;/*MOV    $9  $31  0 */
posHD[994] = 32'b01010111111000000000000000000000;/*OUT    $31  0  */
posHD[995] = 32'b00111000000000000000000000000000;/*JMPR   $0   0  */
posHD[996] = 32'b00110100000000000000001111111001; /*JMP     1017 */
posHD[997] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[998] = 32'b00101000100111100000000000000000;/*MOV    $4  $30  0 */
posHD[999] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[1000] = 32'b00101011110001000000000000000000;/*MOV    $30 $4   0 */
posHD[1001] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[1002] = 32'b00101000100111100000000000000000;/*MOV    $4  $30  0 */
posHD[1003] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[1004] = 32'b00101011110001010000000000000000;/*MOV    $30 $5   0 */
posHD[1005] = 32'b00101000100001000000000000000000;/*MOV    $4  $4   0 */
posHD[1006] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[1007] = 32'b00101011111001010000000000000000;/*MOV    $31 $5   0 */
posHD[1008] = 32'b00101000101001010000000000000000;/*MOV    $5  $5   0 */
posHD[1009] = 32'b01101000000000000000001111101010; /*JAL     1002 */
posHD[1010] = 32'b00101000000111110000000000000000;/*MOV    $0  $31  0 */
posHD[1011] = 32'b10100000000000000000000000000000; /*interrupCPC     0  */

//potencia
posHD[1040] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[1041] = 32'b00110100000000000000010000000011; /*JMP    $1027*/
posHD[1042] = 32'b00100101010000000000000000000001;/*LOI    $10  1  */
posHD[1043] = 32'b00101000000111100000000000000000;/*MOV    $0  $30  0 */
posHD[1044] = 32'b00101000100111100000000000000000;/*MOV    $4  $30  0 */
posHD[1045] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[1046] = 32'b00101001010100010000000000000000;/*MOV    $10 $17  0 */
posHD[1047] = 32'b00101000101111010000000000000000;/*MOV    $5  $29  0 */
posHD[1048] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[1049] = 32'b01001011110111011110100000000000; /*SLET   $30 $29  $29*/
posHD[1050] = 32'b00100111110000000000000000000001;/*LOI    $30  1  */
posHD[1051] = 32'b01000011110111010000001111111111;/*BNEQ   $30 $29  1023*/
posHD[1052] = 32'b00101001001100010000000000000000;/*MOV    $9  $17  0 */
posHD[1053] = 32'b00101000100111010000000000000000;/*MOV    $4  $29  0 */
posHD[1054] = 32'b00101010001111100000000000000000;/*MOV    $17 $30  0 */
posHD[1055] = 32'b01100011101111101111000000000000; /*MULT   $29 $30  $30*/
posHD[1056] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[1057] = 32'b00101011110010010000000000000000;/*MOV    $30 $9   0 */
posHD[1058] = 32'b00101001010100010000000000000000;/*MOV    $10 $17  0 */
posHD[1059] = 32'b00101010001111010000000000000000;/*MOV    $17 $29  0 */
posHD[1060] = 32'b00001011101111100000000000000001;/*ADCI   $29 $30  1 */
posHD[1061] = 32'b00101011110010100000000000000000;/*MOV    $30 $10  0 */
posHD[1062] = 32'b00110100000000000000001111101110; /*JMP     1006 */
posHD[1063] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[1064] = 32'b01011000000000000000000000000000; /*NOP     0  */
posHD[1065] = 32'b00101001001000010000000000000000;/*MOV    $9  $1   0 */
posHD[1066] = 32'b00111000000000000000000000000000;/*JMPR   $0   0  */
posHD[1067] = 32'b00110100000000000000010000000100; /*JMP     1028 */
posHD[1068] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[1069] = 32'b00101000100111100000000000000000;/*MOV    $4  $30  0 */
posHD[1070] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[1071] = 32'b00101011110001000000000000000000;/*MOV    $30 $4   0 */
posHD[1072] = 32'b01010011111000000000000000000000;/*IN     $31  0  */
posHD[1073] = 32'b00101000100111100000000000000000;/*MOV    $4  $30  0 */
posHD[1074] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[1075] = 32'b00101011110001010000000000000000;/*MOV    $30 $5   0 */
posHD[1076] = 32'b00101000100111110000000000000000;/*MOV    $4  $31  0 */
posHD[1077] = 32'b00101000100001000000000000000000;/*MOV    $4  $4   0 */
posHD[1078] = 32'b00101011111111100000000000000000;/*MOV    $31 $30  0 */
posHD[1079] = 32'b00101000101111110000000000000000;/*MOV    $5  $31  0 */
posHD[1080] = 32'b00101011111001010000000000000000;/*MOV    $31 $5   0 */
posHD[1081] = 32'b00101000101001010000000000000000;/*MOV    $5  $5   0 */
posHD[1082] = 32'b01101000000000000000001111101010; /*JAL     1002 */
posHD[1083] = 32'b00101000001111110000000000000000;/*MOV    $1  $31  0 */
posHD[1084] = 32'b01010111111000000000000000000000;/*OUT    $31  0  */
posHD[1085] = 32'b10100000000000000000000000000000; /*interrupCPC     0  */



//retorno do SO

posHD[1100] = 32'b00110100000000000000000000100010; /*JMP     34 */
posHD[1101] = 32'b00110100000000000000000111000100; /*JMP     452 */


end 
	always @ (posedge clk) begin

		if (ONescrita)
				posHD[endereco] = dadoEscrita;
	end
	
	always @ (posedge ck) begin

		dadoLeitura = posHD[endereco];
	end


	
	

endmodule
