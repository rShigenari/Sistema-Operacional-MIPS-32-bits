module UC (opcode, onWriteReg,  writeDataMem, outputEnable, onop, onskip, muxEnd,
ctrlM5, selectSize, selectDado, selectD, HLT, endPCorReg, inputEnable, outmuxReg2,write_mem_inst, save_hd,
reset_pc, writeProcBuffer, flag_inst_type, zerarPC, flagCmd, emit, regType, selectRegFRST, selectReg, onWriteBuf, interrupt);
input [5:0] opcode;
output reg onWriteReg, writeDataMem, outputEnable, onop, onskip, muxEnd, outmuxReg2;
output reg [1:0] ctrlM5, selectSize;
output reg [2:0] selectDado;
output reg selectD, HLT, endPCorReg, inputEnable, write_mem_inst,save_hd, reset_pc, writeProcBuffer ;
output reg [1:0] flag_inst_type;
output reg zerarPC, onWriteBuf; //zerar um pc auxiliar - quantum
output reg flagCmd, emit, regType, selectRegFRST, selectReg, interrupt;

parameter adc = 6'b0, sub = 6'b1, adci = 6'b10, subi = 6'b00011, storePage = 6'b100, loadPage = 6'b101, countPC = 6'b110,
lowo = 6'b00111, stwo = 6'b01000, loi = 6'b1001, mov = 6'b01010, insereInst = 6'b01011, sril = 6'b1100, jump = 6'b1101,
jmpr = 6'b01110, saveProc = 6'b01111, bneq = 6'b10000, blz = 6'b10001, slet = 6'b10010, sgrt = 6'b10011, in = 6'b10100,
out = 6'b10101, nop = 6'b10110, hlt = 6'b10111, mult = 6'b11000, multi = 6'b11001, jal = 6'b11010, div = 6'b11011,
copy = 6'b11100, storeRegister = 6'b011110 , loadRegister = 6'b011101, reset = 6'b11111, inCMD = 6'b100000, emitCMD = 6'b100001,
loi6bits = 6'b100010, savePC = 6'b100011, saveadd_buffer = 6'b100100, renameProg = 6'b100101, troca_contexto = 6'b100110, 
renameProgReg = 6'b100111, interrupCPC  = 6'b101000;

always @ (opcode) begin
	case (opcode)
		adc: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			outmuxReg2 = 0;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			selectDado = 0;
			selectD = 0;
			inputEnable = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;
			onWriteBuf = 0;
			interrupt = 0;
		end
		sub:  begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			outmuxReg2 = 0;
			onop = 1;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			selectDado = 0;
			inputEnable = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;
			onWriteBuf = 0;
			interrupt = 0;
			
		end
		adci:  begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			outmuxReg2 = 0;
			muxEnd = 1;
			inputEnable = 0;
			ctrlM5 = 2'b01;
			selectSize = 2'b0;
			selectDado = 0;
			selectD = 1;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;
			onWriteBuf = 0;
			interrupt = 0;
		end
		subi:
		begin
			onWriteReg = 1;
			writeDataMem = 0;
			inputEnable = 0;
			outputEnable = 0;
			onop = 1;
			outmuxReg2 = 0;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 2'b01;
			selectSize = 2'b0;
			selectDado = 0;
			selectD = 1;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;
			onWriteBuf = 0;
			interrupt = 0;
		end
		storePage: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			outmuxReg2 = 0;
			muxEnd = 1;
			ctrlM5 = 2'b10;
			inputEnable = 0;
			selectSize = 2'bx;
			selectDado = 0;
			selectD = 0;	
			writeProcBuffer = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;
			onWriteBuf = 0;
			interrupt = 0;
		end
		loadPage:  begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			inputEnable = 0;
			outmuxReg2 = 0;
			muxEnd = 1;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b10;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;		
		   onWriteBuf = 0;	
			interrupt = 0;
		end
	countPC: begin //na troca de contexto, lançar instrucao de countPC e fazer jr
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			outmuxReg2 = 0;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 2'b01;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 1;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		
	lowo: begin
			writeProcBuffer = 0;
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			inputEnable = 0;
			outmuxReg2 = 1;
			muxEnd = 1;
			ctrlM5 = 2'b10;
			selectSize = 2'b0;
			selectDado = 3'b10;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		stwo: begin
			onWriteReg = 0;
			writeDataMem = 1;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			outmuxReg2 = 1;
			inputEnable = 0;
			muxEnd = 1;
			ctrlM5 = 2'bx;
			selectSize = 2'b0;
			selectDado = 2'bx;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		loi: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			outmuxReg2 = 0;
			inputEnable = 0;
			muxEnd = 1;
			ctrlM5 = 0;
			selectSize = 2'b01;
			selectDado = 3'b11;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		mov: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			outmuxReg2 = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			inputEnable = 0;
			ctrlM5 = 2'b01;
			selectSize = 2'bx;
			selectDado = 3'b01;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		insereInst: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			outmuxReg2 = 0;
			muxEnd = 1;
			ctrlM5 = 2'b01;
			inputEnable = 0;
			selectSize = 2'b0;
			selectDado = 0;
			selectD = 1;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		sril: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			muxEnd = 1;
			inputEnable = 0;
			outmuxReg2 = 0;
			ctrlM5 = 1;
			selectSize = 2'b0;
			selectDado = 0;
			selectD = 1;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		jump: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			outmuxReg2 = 0;
			inputEnable = 0;
			onop = 0;
			onskip = 1;
			muxEnd = 0;
			ctrlM5 = 2'bx;
			selectSize = 2'bx;
			selectDado = 3'bx;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		jmpr: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 1;
			muxEnd = 0;
			outmuxReg2 = 0;
			ctrlM5 = 0;
			selectSize = 0;
			selectDado = 0;
			selectD = 0;
			inputEnable = 0;
			HLT = 0;
			endPCorReg = 1;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		saveProc: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			outmuxReg2 = 0;
			onskip = 0;
			muxEnd = 0;
			ctrlM5 = 2'bx;
			inputEnable = 0;
			selectSize = 2'bx;
			selectDado = 2'bx;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 1;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		bneq: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			outmuxReg2 = 0;
			onop = 1;
			onskip = 1;
			muxEnd = 0;
			ctrlM5 = 2'bx;
			inputEnable = 0;
			selectSize = 2'bx;
			selectDado = 2'bx;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		blz: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			outmuxReg2 = 0;
			inputEnable = 0;
			onskip = 1;
			muxEnd = 0;
			ctrlM5 = 2'bx;
			selectSize = 2'bx;
			selectDado = 2'bx;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		slet: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			inputEnable = 0;
			outmuxReg2 = 0;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		sgrt: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			inputEnable = 0;
			onskip = 0;
			outmuxReg2 = 0;
			muxEnd = 1;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		in: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			inputEnable = 1;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b0;
			selectSize = 2'b11;
			selectDado = 3'b11;
			selectD = 1;
			HLT = 1;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		out: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 1;
			outmuxReg2 = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 2'bx;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 3'bx;
			selectD = 1'bx;
			HLT = 1;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		nop:
		begin
			onWriteReg = 0;
			writeDataMem = 0;
			inputEnable = 0;
			outmuxReg2 = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 0;
			selectSize = 2'b0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		hlt: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			outmuxReg2 = 0;
			onskip = 0;
			muxEnd = 1;
			inputEnable = 0;
			ctrlM5 = 2'bx;
			selectSize = 2'bx;
			selectDado = 2'bx;
			selectD = 1'bx;
			HLT = 1;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		mult: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
			multi: begin
			onWriteReg = 1;
			writeDataMem = 0;
			inputEnable = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			muxEnd = 1;
			ctrlM5 = 2'b01;
			outmuxReg2 = 0;
			selectSize = 2'b0;
			selectDado = 0;
			selectD = 1;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 3'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
			end

			jal: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 1;
			muxEnd = 0;
			ctrlM5 = 2'b00;
			selectSize = 2'b10;
			outmuxReg2 = 0;
			inputEnable = 0;
			selectDado = 3'b11;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end

		div: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 1;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end

		copy: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 1;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b0;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end

		storeRegister: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 1;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b1;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 1;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		
		loadRegister: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b11;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 3'b100;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b1;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 1;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		
		reset: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 1;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		inCMD: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'b11;
			inputEnable = 1;
			selectDado = 3'b11;
			selectD = 1;
			HLT = 1;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 1;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		emitCMD: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 1;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		
		loi6bits: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			outmuxReg2 = 0;
			inputEnable = 0;
			muxEnd = 1;
			ctrlM5 = 0;
			selectSize = 2'b0;
			selectDado = 3'b11;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 1;
			emit = 0;
			regType = 1;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		
		renameProgReg: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			outmuxReg2 = 0;
			inputEnable = 0;
			muxEnd = 1;
			ctrlM5 = 0;
			selectSize = 2'b0;
			selectDado = 3'b11;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 1;
			interrupt = 0;
		end 
		
		troca_contexto: begin
			onWriteReg = 1;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			outmuxReg2 = 0;
			inputEnable = 0;
			muxEnd = 1;
			ctrlM5 = 2'b1;
			selectSize = 2'b0;
			selectDado = 3'b101;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
			
		end 
		
		interrupCPC: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			outmuxReg2 = 0;
			inputEnable = 0;
			muxEnd = 1;
			ctrlM5 = 2'b1;
			selectSize = 2'b0;
			selectDado = 3'b101;
			selectD = 1'bx;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 1;
			
		end 
		


		default: begin
			onWriteReg = 0;
			writeDataMem = 0;
			outputEnable = 0;
			onop = 0;
			onskip = 0;
			muxEnd = 1;
			outmuxReg2 = 0;
			ctrlM5 = 2'b10;
			selectSize = 2'bx;
			inputEnable = 0;
			selectDado = 0;
			selectD = 0;
			HLT = 0;
			endPCorReg = 0;
			write_mem_inst= 0;
			save_hd = 0;
			reset_pc = 0;
			writeProcBuffer = 0;
			flag_inst_type = 2'b11;
			zerarPC = 0;
			flagCmd = 0;
			emit = 0;
			regType = 0;
			selectRegFRST = 0;
			selectReg = 0;	
			onWriteBuf = 0;
			interrupt = 0;
		end
		
	
	endcase
end

endmodule
